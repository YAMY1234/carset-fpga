`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2020/12/28 08:52:55
// Design Name: 
// Module Name: read_bg_data
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


/*
$fseek���ļ���λ�����Դ��������ļ����в�����

$fscanf�����ļ�һ�н��ж�д��
*/


module read_bg_data(
    
    );
endmodule
